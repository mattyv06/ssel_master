.title KiCad schematic
.include "LTC1044A.sub"
.include "sub/diode/sdm10m45sd.sub"
.include "sub/sim/beh_iload.sub"
Vin1 /CHARGE_PUMP/PWR_IN 0 dc 6
Ictl1 0 /L1 dc 10m
XB1 /CHARGE_PUMP/PWR_OUT /L1 beh_iload
CC2 /CHARGE_PUMP/D1 /CHARGE_PUMP/CAP 10u
CC3 /CHARGE_PUMP/D2 0 10u
CC1 /CHARGE_PUMP/PWR_IN 0 100n
XU1 nc1 /CHARGE_PUMP/CAP 0 nc2 nc3 nc4 nc5 /CHARGE_PUMP/PWR_IN LTC1044A
CC4 /CHARGE_PUMP/D3 /CHARGE_PUMP/CAP 10u
CC5 /CHARGE_PUMP/PWR_OUT 0 10u
XD1 /CHARGE_PUMP/PWR_IN /CHARGE_PUMP/D2 /CHARGE_PUMP/D3 /CHARGE_PUMP/D2 /CHARGE_PUMP/PWR_OUT /CHARGE_PUMP/D1 SDM10M45SD
.tran 100m
.step Vin1 5.5 8.5 1
.end
